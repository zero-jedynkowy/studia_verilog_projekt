module exe_unit_w1(i_oper, i_argA, i_argB, i_clk, i_rsn, o_result, o_status);
    input logic [n:0] i_oper;
    input logic [m:0] i_argA;
    input logic [m:0] i_argB;
    input logic i_clk;
    input logic i_rsn;
    output logic [m:0] o_result;
    output logic [2:0] o_status;
    //test
endmodule